component mosquitto.Printnum

endpoints {
    printnum : mosquitto.Printnum
}